/*
 * A simple fake RAM that you can use to aid in debugging your wave display.
 */
module fake_sample_ram (
    input clk,
    input [8:0] addr,
    output reg [7:0] dout
);

    always @(posedge clk)
            dout = memory[addr];
    

	wire [7:0] memory [511:0];			
	assign memory[	  0	] =	8'd128;
	assign memory[	  1	] =	8'd141;
	assign memory[	  2	] =	8'd153;
	assign memory[	  3	] =	8'd166;
	assign memory[	  4	] =	8'd177;
	assign memory[	  5	] =	8'd189;
	assign memory[	  6	] =	8'd200;
	assign memory[	  7	] =	8'd210;
	assign memory[	  8	] =	8'd219;
	assign memory[	  9	] =	8'd227;
	assign memory[	 10	] =	8'd235;
	assign memory[	 11	] =	8'd241;
	assign memory[	 12	] =	8'd246;
	assign memory[	 13	] =	8'd250;
	assign memory[	 14	] =	8'd253;
	assign memory[	 15	] =	8'd255;
	assign memory[	 16	] =	8'd255;
	assign memory[	 17	] =	8'd254;
	assign memory[	 18	] =	8'd252;
	assign memory[	 19	] =	8'd248;
	assign memory[	 20	] =	8'd243;
	assign memory[	 21	] =	8'd238;
	assign memory[	 22	] =	8'd231;
	assign memory[	 23	] =	8'd223;
	assign memory[	 24	] =	8'd214;
	assign memory[	 25	] =	8'd204;
	assign memory[	 26	] =	8'd193;
	assign memory[	 27	] =	8'd182;
	assign memory[	 28	] =	8'd171;
	assign memory[	 29	] =	8'd158;
	assign memory[	 30	] =	8'd146;
	assign memory[	 31	] =	8'd133;
	assign memory[	 32	] =	8'd121;
	assign memory[	 33	] =	8'd108;
	assign memory[	 34	] =	8'd96;
	assign memory[	 35	] =	8'd83;
	assign memory[	 36	] =	8'd72;
	assign memory[	 37	] =	8'd61;
	assign memory[	 38	] =	8'd50;
	assign memory[	 39	] =	8'd41;
	assign memory[	 40	] =	8'd32;
	assign memory[	 41	] =	8'd24;
	assign memory[	 42	] =	8'd17;
	assign memory[	 43	] =	8'd12;
	assign memory[	 44	] =	8'd7;
	assign memory[	 45	] =	8'd4;
	assign memory[	 46	] =	8'd2;
	assign memory[	 47	] =	8'd1;
	assign memory[	 48	] =	8'd1;
	assign memory[	 49	] =	8'd3;
	assign memory[	 50	] =	8'd6;
	assign memory[	 51	] =	8'd10;
	assign memory[	 52	] =	8'd16;
	assign memory[	 53	] =	8'd22;
	assign memory[	 54	] =	8'd30;
	assign memory[	 55	] =	8'd38;
	assign memory[	 56	] =	8'd48;
	assign memory[	 57	] =	8'd58;
	assign memory[	 58	] =	8'd69;
	assign memory[	 59	] =	8'd81;
	assign memory[	 60	] =	8'd93;
	assign memory[	 61	] =	8'd105;
	assign memory[	 62	] =	8'd117;
	assign memory[	 63	] =	8'd130;
	assign memory[	 64	] =	8'd143;
	assign memory[	 65	] =	8'd155;
	assign memory[	 66	] =	8'd168;
	assign memory[	 67	] =	8'd179;
	assign memory[	 68	] =	8'd191;
	assign memory[	 69	] =	8'd201;
	assign memory[	 70	] =	8'd211;
	assign memory[	 71	] =	8'd221;
	assign memory[	 72	] =	8'd229;
	assign memory[	 73	] =	8'd236;
	assign memory[	 74	] =	8'd242;
	assign memory[	 75	] =	8'd247;
	assign memory[	 76	] =	8'd251;
	assign memory[	 77	] =	8'd253;
	assign memory[	 78	] =	8'd255;
	assign memory[	 79	] =	8'd255;
	assign memory[	 80	] =	8'd254;
	assign memory[	 81	] =	8'd251;
	assign memory[	 82	] =	8'd247;
	assign memory[	 83	] =	8'd243;
	assign memory[	 84	] =	8'd237;
	assign memory[	 85	] =	8'd229;
	assign memory[	 86	] =	8'd221;
	assign memory[	 87	] =	8'd212;
	assign memory[	 88	] =	8'd202;
	assign memory[	 89	] =	8'd192;
	assign memory[	 90	] =	8'd180;
	assign memory[	 91	] =	8'd169;
	assign memory[	 92	] =	8'd156;
	assign memory[	 93	] =	8'd144;
	assign memory[	 94	] =	8'd131;
	assign memory[	 95	] =	8'd118;
	assign memory[	 96	] =	8'd106;
	assign memory[	 97	] =	8'd93;
	assign memory[	 98	] =	8'd81;
	assign memory[	 99	] =	8'd70;
	assign memory[	100	] =	8'd59;
	assign memory[	101	] =	8'd49;
	assign memory[	102	] =	8'd39;
	assign memory[	103	] =	8'd31;
	assign memory[	104	] =	8'd23;
	assign memory[	105	] =	8'd16;
	assign memory[	106	] =	8'd11;
	assign memory[	107	] =	8'd7;
	assign memory[	108	] =	8'd3;
	assign memory[	109	] =	8'd2;
	assign memory[	110	] =	8'd1;
	assign memory[	111	] =	8'd2;
	assign memory[	112	] =	8'd4;
	assign memory[	113	] =	8'd7;
	assign memory[	114	] =	8'd11;
	assign memory[	115	] =	8'd17;
	assign memory[	116	] =	8'd24;
	assign memory[	117	] =	8'd31;
	assign memory[	118	] =	8'd40;
	assign memory[	119	] =	8'd49;
	assign memory[	120	] =	8'd60;
	assign memory[	121	] =	8'd71;
	assign memory[	122	] =	8'd83;
	assign memory[	123	] =	8'd95;
	assign memory[	124	] =	8'd107;
	assign memory[	125	] =	8'd120;
	assign memory[	126	] =	8'd132;
	assign memory[	127	] =	8'd145;
	assign memory[	128	] =	8'd157;
	assign memory[	129	] =	8'd170;
	assign memory[	130	] =	8'd181;
	assign memory[	131	] =	8'd193;
	assign memory[	132	] =	8'd203;
	assign memory[	133	] =	8'd213;
	assign memory[	134	] =	8'd222;
	assign memory[	135	] =	8'd230;
	assign memory[	136	] =	8'd237;
	assign memory[	137	] =	8'd243;
	assign memory[	138	] =	8'd248;
	assign memory[	139	] =	8'd251;
	assign memory[	140	] =	8'd254;
	assign memory[	141	] =	8'd255;
	assign memory[	142	] =	8'd255;
	assign memory[	143	] =	8'd253;
	assign memory[	144	] =	8'd251;
	assign memory[	145	] =	8'd247;
	assign memory[	146	] =	8'd242;
	assign memory[	147	] =	8'd235;
	assign memory[	148	] =	8'd228;
	assign memory[	149	] =	8'd220;
	assign memory[	150	] =	8'd211;
	assign memory[	151	] =	8'd201;
	assign memory[	152	] =	8'd190;
	assign memory[	153	] =	8'd178;
	assign memory[	154	] =	8'd166;
	assign memory[	155	] =	8'd154;
	assign memory[	156	] =	8'd142;
	assign memory[	157	] =	8'd129;
	assign memory[	158	] =	8'd116;
	assign memory[	159	] =	8'd104;
	assign memory[	160	] =	8'd91;
	assign memory[	161	] =	8'd79;
	assign memory[	162	] =	8'd68;
	assign memory[	163	] =	8'd57;
	assign memory[	164	] =	8'd47;
	assign memory[	165	] =	8'd38;
	assign memory[	166	] =	8'd29;
	assign memory[	167	] =	8'd22;
	assign memory[	168	] =	8'd15;
	assign memory[	169	] =	8'd10;
	assign memory[	170	] =	8'd6;
	assign memory[	171	] =	8'd3;
	assign memory[	172	] =	8'd1;
	assign memory[	173	] =	8'd1;
	assign memory[	174	] =	8'd2;
	assign memory[	175	] =	8'd4;
	assign memory[	176	] =	8'd7;
	assign memory[	177	] =	8'd12;
	assign memory[	178	] =	8'd18;
	assign memory[	179	] =	8'd25;
	assign memory[	180	] =	8'd33;
	assign memory[	181	] =	8'd41;
	assign memory[	182	] =	8'd51;
	assign memory[	183	] =	8'd62;
	assign memory[	184	] =	8'd73;
	assign memory[	185	] =	8'd85;
	assign memory[	186	] =	8'd97;
	assign memory[	187	] =	8'd109;
	assign memory[	188	] =	8'd122;
	assign memory[	189	] =	8'd134;
	assign memory[	190	] =	8'd147;
	assign memory[	191	] =	8'd159;
	assign memory[	192	] =	8'd172;
	assign memory[	193	] =	8'd183;
	assign memory[	194	] =	8'd194;
	assign memory[	195	] =	8'd205;
	assign memory[	196	] =	8'd215;
	assign memory[	197	] =	8'd223;
	assign memory[	198	] =	8'd231;
	assign memory[	199	] =	8'd238;
	assign memory[	200	] =	8'd244;
	assign memory[	201	] =	8'd249;
	assign memory[	202	] =	8'd252;
	assign memory[	203	] =	8'd254;
	assign memory[	204	] =	8'd255;
	assign memory[	205	] =	8'd255;
	assign memory[	206	] =	8'd253;
	assign memory[	207	] =	8'd250;
	assign memory[	208	] =	8'd246;
	assign memory[	209	] =	8'd241;
	assign memory[	210	] =	8'd234;
	assign memory[	211	] =	8'd227;
	assign memory[	212	] =	8'd218;
	assign memory[	213	] =	8'd209;
	assign memory[	214	] =	8'd199;
	assign memory[	215	] =	8'd188;
	assign memory[	216	] =	8'd176;
	assign memory[	217	] =	8'd164;
	assign memory[	218	] =	8'd152;
	assign memory[	219	] =	8'd140;
	assign memory[	220	] =	8'd127;
	assign memory[	221	] =	8'd114;
	assign memory[	222	] =	8'd102;
	assign memory[	223	] =	8'd89;
	assign memory[	224	] =	8'd78;
	assign memory[	225	] =	8'd66;
	assign memory[	226	] =	8'd55;
	assign memory[	227	] =	8'd45;
	assign memory[	228	] =	8'd36;
	assign memory[	229	] =	8'd28;
	assign memory[	230	] =	8'd21;
	assign memory[	231	] =	8'd14;
	assign memory[	232	] =	8'd9;
	assign memory[	233	] =	8'd5;
	assign memory[	234	] =	8'd3;
	assign memory[	235	] =	8'd1;
	assign memory[	236	] =	8'd1;
	assign memory[	237	] =	8'd2;
	assign memory[	238	] =	8'd5;
	assign memory[	239	] =	8'd8;
	assign memory[	240	] =	8'd13;
	assign memory[	241	] =	8'd19;
	assign memory[	242	] =	8'd26;
	assign memory[	243	] =	8'd34;
	assign memory[	244	] =	8'd43;
	assign memory[	245	] =	8'd53;
	assign memory[	246	] =	8'd63;
	assign memory[	247	] =	8'd75;
	assign memory[	248	] =	8'd87;
	assign memory[	249	] =	8'd99;
	assign memory[	250	] =	8'd111;
	assign memory[	251	] =	8'd124;
	assign memory[	252	] =	8'd137;
	assign memory[	253	] =	8'd149;
	assign memory[	254	] =	8'd162;
	assign memory[	255	] =	8'd174;
	assign memory[	256	] =	8'd185;
	assign memory[	257	] =	8'd196;
	assign memory[	258	] =	8'd207;
	assign memory[	259	] =	8'd216;
	assign memory[	260	] =	8'd225;
	assign memory[	261	] =	8'd233;
	assign memory[	262	] =	8'd239;
	assign memory[	263	] =	8'd245;
	assign memory[	264	] =	8'd249;
	assign memory[	265	] =	8'd252;
	assign memory[	266	] =	8'd254;
	assign memory[	267	] =	8'd255;
	assign memory[	268	] =	8'd254;
	assign memory[	269	] =	8'd253;
	assign memory[	270	] =	8'd249;
	assign memory[	271	] =	8'd245;
	assign memory[	272	] =	8'd240;
	assign memory[	273	] =	8'd233;
	assign memory[	274	] =	8'd225;
	assign memory[	275	] =	8'd217;
	assign memory[	276	] =	8'd207;
	assign memory[	277	] =	8'd197;
	assign memory[	278	] =	8'd186;
	assign memory[	279	] =	8'd174;
	assign memory[	280	] =	8'd162;
	assign memory[	281	] =	8'd150;
	assign memory[	282	] =	8'd137;
	assign memory[	283	] =	8'd125;
	assign memory[	284	] =	8'd112;
	assign memory[	285	] =	8'd100;
	assign memory[	286	] =	8'd87;
	assign memory[	287	] =	8'd76;
	assign memory[	288	] =	8'd64;
	assign memory[	289	] =	8'd54;
	assign memory[	290	] =	8'd44;
	assign memory[	291	] =	8'd35;
	assign memory[	292	] =	8'd27;
	assign memory[	293	] =	8'd19;
	assign memory[	294	] =	8'd13;
	assign memory[	295	] =	8'd8;
	assign memory[	296	] =	8'd5;
	assign memory[	297	] =	8'd2;
	assign memory[	298	] =	8'd1;
	assign memory[	299	] =	8'd1;
	assign memory[	300	] =	8'd3;
	assign memory[	301	] =	8'd5;
	assign memory[	302	] =	8'd9;
	assign memory[	303	] =	8'd14;
	assign memory[	304	] =	8'd20;
	assign memory[	305	] =	8'd27;
	assign memory[	306	] =	8'd35;
	assign memory[	307	] =	8'd45;
	assign memory[	308	] =	8'd55;
	assign memory[	309	] =	8'd65;
	assign memory[	310	] =	8'd77;
	assign memory[	311	] =	8'd89;
	assign memory[	312	] =	8'd101;
	assign memory[	313	] =	8'd113;
	assign memory[	314	] =	8'd126;
	assign memory[	315	] =	8'd139;
	assign memory[	316	] =	8'd151;
	assign memory[	317	] =	8'd164;
	assign memory[	318	] =	8'd176;
	assign memory[	319	] =	8'd187;
	assign memory[	320	] =	8'd198;
	assign memory[	321	] =	8'd208;
	assign memory[	322	] =	8'd218;
	assign memory[	323	] =	8'd226;
	assign memory[	324	] =	8'd234;
	assign memory[	325	] =	8'd240;
	assign memory[	326	] =	8'd246;
	assign memory[	327	] =	8'd250;
	assign memory[	328	] =	8'd253;
	assign memory[	329	] =	8'd255;
	assign memory[	330	] =	8'd255;
	assign memory[	331	] =	8'd254;
	assign memory[	332	] =	8'd252;
	assign memory[	333	] =	8'd249;
	assign memory[	334	] =	8'd244;
	assign memory[	335	] =	8'd239;
	assign memory[	336	] =	8'd232;
	assign memory[	337	] =	8'd224;
	assign memory[	338	] =	8'd215;
	assign memory[	339	] =	8'd206;
	assign memory[	340	] =	8'd195;
	assign memory[	341	] =	8'd184;
	assign memory[	342	] =	8'd172;
	assign memory[	343	] =	8'd160;
	assign memory[	344	] =	8'd148;
	assign memory[	345	] =	8'd135;
	assign memory[	346	] =	8'd123;
	assign memory[	347	] =	8'd110;
	assign memory[	348	] =	8'd98;
	assign memory[	349	] =	8'd85;
	assign memory[	350	] =	8'd74;
	assign memory[	351	] =	8'd62;
	assign memory[	352	] =	8'd52;
	assign memory[	353	] =	8'd42;
	assign memory[	354	] =	8'd33;
	assign memory[	355	] =	8'd25;
	assign memory[	356	] =	8'd18;
	assign memory[	357	] =	8'd12;
	assign memory[	358	] =	8'd8;
	assign memory[	359	] =	8'd4;
	assign memory[	360	] =	8'd2;
	assign memory[	361	] =	8'd1;
	assign memory[	362	] =	8'd1;
	assign memory[	363	] =	8'd3;
	assign memory[	364	] =	8'd6;
	assign memory[	365	] =	8'd10;
	assign memory[	366	] =	8'd15;
	assign memory[	367	] =	8'd21;
	assign memory[	368	] =	8'd29;
	assign memory[	369	] =	8'd37;
	assign memory[	370	] =	8'd46;
	assign memory[	371	] =	8'd56;
	assign memory[	372	] =	8'd67;
	assign memory[	373	] =	8'd79;
	assign memory[	374	] =	8'd91;
	assign memory[	375	] =	8'd103;
	assign memory[	376	] =	8'd115;
	assign memory[	377	] =	8'd128;
	assign memory[	378	] =	8'd141;
	assign memory[	379	] =	8'd153;
	assign memory[	380	] =	8'd166;
	assign memory[	381	] =	8'd178;
	assign memory[	382	] =	8'd189;
	assign memory[	383	] =	8'd200;
	assign memory[	384	] =	8'd210;
	assign memory[	385	] =	8'd219;
	assign memory[	386	] =	8'd228;
	assign memory[	387	] =	8'd235;
	assign memory[	388	] =	8'd241;
	assign memory[	389	] =	8'd246;
	assign memory[	390	] =	8'd250;
	assign memory[	391	] =	8'd253;
	assign memory[	392	] =	8'd255;
	assign memory[	393	] =	8'd255;
	assign memory[	394	] =	8'd254;
	assign memory[	395	] =	8'd252;
	assign memory[	396	] =	8'd248;
	assign memory[	397	] =	8'd243;
	assign memory[	398	] =	8'd238;
	assign memory[	399	] =	8'd231;
	assign memory[	400	] =	8'd223;
	assign memory[	401	] =	8'd214;
	assign memory[	402	] =	8'd204;
	assign memory[	403	] =	8'd193;
	assign memory[	404	] =	8'd182;
	assign memory[	405	] =	8'd170;
	assign memory[	406	] =	8'd158;
	assign memory[	407	] =	8'd146;
	assign memory[	408	] =	8'd133;
	assign memory[	409	] =	8'd120;
	assign memory[	410	] =	8'd108;
	assign memory[	411	] =	8'd95;
	assign memory[	412	] =	8'd83;
	assign memory[	413	] =	8'd72;
	assign memory[	414	] =	8'd61;
	assign memory[	415	] =	8'd50;
	assign memory[	416	] =	8'd41;
	assign memory[	417	] =	8'd32;
	assign memory[	418	] =	8'd24;
	assign memory[	419	] =	8'd17;
	assign memory[	420	] =	8'd12;
	assign memory[	421	] =	8'd7;
	assign memory[	422	] =	8'd4;
	assign memory[	423	] =	8'd2;
	assign memory[	424	] =	8'd1;
	assign memory[	425	] =	8'd1;
	assign memory[	426	] =	8'd3;
	assign memory[	427	] =	8'd6;
	assign memory[	428	] =	8'd10;
	assign memory[	429	] =	8'd16;
	assign memory[	430	] =	8'd22;
	assign memory[	431	] =	8'd30;
	assign memory[	432	] =	8'd38;
	assign memory[	433	] =	8'd48;
	assign memory[	434	] =	8'd58;
	assign memory[	435	] =	8'd69;
	assign memory[	436	] =	8'd81;
	assign memory[	437	] =	8'd93;
	assign memory[	438	] =	8'd105;
	assign memory[	439	] =	8'd118;
	assign memory[	440	] =	8'd130;
	assign memory[	441	] =	8'd143;
	assign memory[	442	] =	8'd155;
	assign memory[	443	] =	8'd168;
	assign memory[	444	] =	8'd180;
	assign memory[	445	] =	8'd191;
	assign memory[	446	] =	8'd202;
	assign memory[	447	] =	8'd212;
	assign memory[	448	] =	8'd221;
	assign memory[	449	] =	8'd229;
	assign memory[	450	] =	8'd236;
	assign memory[	451	] =	8'd242;
	assign memory[	452	] =	8'd247;
	assign memory[	453	] =	8'd251;
	assign memory[	454	] =	8'd254;
	assign memory[	455	] =	8'd255;
	assign memory[	456	] =	8'd255;
	assign memory[	457	] =	8'd254;
	assign memory[	458	] =	8'd251;
	assign memory[	459	] =	8'd247;
	assign memory[	460	] =	8'd243;
	assign memory[	461	] =	8'd236;
	assign memory[	462	] =	8'd229;
	assign memory[	463	] =	8'd221;
	assign memory[	464	] =	8'd212;
	assign memory[	465	] =	8'd202;
	assign memory[	466	] =	8'd192;
	assign memory[	467	] =	8'd180;
	assign memory[	468	] =	8'd168;
	assign memory[	469	] =	8'd156;
	assign memory[	470	] =	8'd144;
	assign memory[	471	] =	8'd131;
	assign memory[	472	] =	8'd118;
	assign memory[	473	] =	8'd106;
	assign memory[	474	] =	8'd93;
	assign memory[	475	] =	8'd81;
	assign memory[	476	] =	8'd70;
	assign memory[	477	] =	8'd59;
	assign memory[	478	] =	8'd49;
	assign memory[	479	] =	8'd39;
	assign memory[	480	] =	8'd30;
	assign memory[	481	] =	8'd23;
	assign memory[	482	] =	8'd16;
	assign memory[	483	] =	8'd11;
	assign memory[	484	] =	8'd6;
	assign memory[	485	] =	8'd3;
	assign memory[	486	] =	8'd2;
	assign memory[	487	] =	8'd1;
	assign memory[	488	] =	8'd2;
	assign memory[	489	] =	8'd4;
	assign memory[	490	] =	8'd7;
	assign memory[	491	] =	8'd11;
	assign memory[	492	] =	8'd17;
	assign memory[	493	] =	8'd24;
	assign memory[	494	] =	8'd31;
	assign memory[	495	] =	8'd40;
	assign memory[	496	] =	8'd50;
	assign memory[	497	] =	8'd60;
	assign memory[	498	] =	8'd71;
	assign memory[	499	] =	8'd83;
	assign memory[	500	] =	8'd95;
	assign memory[	501	] =	8'd107;
	assign memory[	502	] =	8'd120;
	assign memory[	503	] =	8'd132;
	assign memory[	504	] =	8'd145;
	assign memory[	505	] =	8'd158;
	assign memory[	506	] =	8'd170;
	assign memory[	507	] =	8'd181;
	assign memory[	508	] =	8'd193;
	assign memory[	509	] =	8'd203;
	assign memory[	510	] =	8'd213;
	assign memory[	511	] =	8'd222;


endmodule				


